module writeback();



endmodule