module sc_logic(next_state, state, rst, err)
	input rst
	input [2:0] state;
	reg [2:0] next_state;
	reg error;
	
endmodule